magic
tech scmos
timestamp 0
use router_generated_wiring gen_wiring
timestamp 976159489
transform 1 0 0 0 1 0
box 0 0 25 61
<< metal1 >>
rect 21 0 24 7
rect 14 0 17 7
rect 7 0 10 7
rect 0 0 3 7
rect 21 56 24 63
rect 14 56 17 63
rect 7 56 10 63
rect 0 56 3 63
<< metal2 >>
rect 21 0 24 7
rect 14 0 17 7
rect 7 0 10 7
rect 0 0 3 7
rect 21 56 24 63
rect 14 56 17 63
rect 7 56 10 63
rect 0 56 3 63
<< labels >>
rlabel metal1 22 58 22 58 1 x7
rlabel metal1 15 60 15 60 3 x5
rlabel metal1 9 60 9 60 3 x3
rlabel metal1 2 59 2 59 3 x1
rlabel metal2 22 59 22 59 7 x8
rlabel metal2 16 58 16 58 1 x6
rlabel metal2 8 60 8 60 3 x4
rlabel metal2 1 60 1 60 3 x2
rlabel metal1 22 2 22 2 1 x7
rlabel metal1 15 4 15 4 3 x5
rlabel metal1 9 4 9 4 3 x3
rlabel metal1 2 3 2 3 3 x1
rlabel metal2 22 3 22 3 7 x8
rlabel metal2 16 2 16 2 1 x6
rlabel metal2 8 4 8 4 3 x4
rlabel metal2 1 4 1 4 3 x2
<< end >>
