magic
tech scmos
timestamp 976159201
<< error_s >>
rect 10 132 11 133
rect 31 132 32 133
rect 54 132 55 133
rect 91 132 92 133
rect 9 131 10 132
rect 32 131 34 132
rect 52 131 54 132
rect 92 131 93 132
rect 34 130 35 131
rect 51 130 52 131
rect 265 130 266 131
rect 286 130 287 131
rect 9 129 10 130
rect 92 129 93 130
rect 264 129 265 130
rect 287 129 289 130
rect 10 128 11 129
rect 91 128 92 129
rect 289 128 290 129
rect 23 127 24 128
rect 62 127 63 128
rect 264 127 265 128
rect 24 126 26 127
rect 60 126 62 127
rect 265 126 266 127
rect 26 125 27 126
rect 59 125 60 126
rect 278 125 279 126
rect 279 124 281 125
rect 281 123 282 124
rect 10 122 11 123
rect 15 122 16 123
rect 86 122 87 123
rect 91 122 92 123
rect 9 121 10 122
rect 16 121 18 122
rect 84 121 86 122
rect 92 121 93 122
rect 18 120 19 121
rect 83 120 84 121
rect 265 120 266 121
rect 270 120 271 121
rect 264 119 265 120
rect 271 119 273 120
rect 273 118 274 119
rect 9 116 10 117
rect 92 116 93 117
rect 10 115 11 116
rect 91 115 92 116
rect 264 114 265 115
rect 265 113 266 114
rect 10 106 11 107
rect 91 106 92 107
rect 9 105 10 106
rect 92 105 93 106
rect 265 104 266 105
rect 264 103 265 104
rect 18 101 19 102
rect 83 101 84 102
rect 9 100 10 101
rect 16 100 18 101
rect 84 100 86 101
rect 92 100 93 101
rect 10 99 11 100
rect 15 99 16 100
rect 86 99 87 100
rect 91 99 92 100
rect 273 99 274 100
rect 264 98 265 99
rect 271 98 273 99
rect 265 97 266 98
rect 270 97 271 98
rect 26 96 27 97
rect 59 96 60 97
rect 24 95 26 96
rect 60 95 62 96
rect 23 94 24 95
rect 62 94 63 95
rect 281 94 282 95
rect 10 93 11 94
rect 91 93 92 94
rect 279 93 281 94
rect 9 92 10 93
rect 92 92 93 93
rect 278 92 279 93
rect 34 91 35 92
rect 51 91 52 92
rect 265 91 266 92
rect 9 90 10 91
rect 32 90 34 91
rect 52 90 54 91
rect 92 90 93 91
rect 264 90 265 91
rect 10 89 11 90
rect 31 89 32 90
rect 54 89 55 90
rect 91 89 92 90
rect 289 89 290 90
rect 264 88 265 89
rect 287 88 289 89
rect 265 87 266 88
rect 286 87 287 88
rect 49 81 57 85
rect 49 77 53 81
rect 31 76 32 77
rect 67 76 68 77
rect 99 76 100 78
rect 32 75 34 76
rect 65 75 67 76
rect 34 74 35 75
rect 64 74 65 75
rect 286 74 287 75
rect 287 73 289 74
rect 2 71 3 73
rect 26 71 27 72
rect 28 71 29 73
rect 72 71 73 72
rect 27 70 29 71
rect 31 70 32 71
rect 70 70 72 71
rect 28 69 30 70
rect 28 68 29 69
rect 2 66 3 68
rect 18 66 19 67
rect 41 66 42 70
rect 69 69 70 70
rect 98 69 102 73
rect 289 72 290 73
rect 257 69 258 71
rect 281 69 282 70
rect 282 68 284 69
rect 284 67 285 68
rect 80 66 81 67
rect 19 65 21 66
rect 78 65 80 66
rect 21 64 22 65
rect 77 64 78 65
rect 257 64 258 66
rect 273 64 274 65
rect 274 63 276 64
rect 13 61 14 62
rect 14 60 16 61
rect 16 59 17 60
rect 41 59 42 63
rect 85 61 86 62
rect 99 61 100 63
rect 276 62 277 63
rect 83 60 85 61
rect 82 59 83 60
rect 39 56 40 59
rect 238 56 242 60
rect 268 59 269 60
rect 269 58 271 59
rect 271 57 272 58
rect 37 53 38 56
rect 41 55 42 56
rect 41 54 45 55
rect 0 49 4 53
rect 25 50 27 51
rect 30 50 31 51
rect 35 50 39 51
rect 41 50 42 54
rect 19 47 20 50
rect 24 48 25 49
rect 27 48 28 50
rect 30 49 39 50
rect 54 49 55 52
rect 56 49 57 51
rect 238 49 242 53
rect 30 48 37 49
rect 280 48 282 49
rect 25 47 26 48
rect 31 46 34 48
rect 0 42 4 46
rect 33 44 34 46
rect 35 44 37 46
rect 22 42 27 43
rect 30 42 32 43
rect 41 42 42 44
rect 238 42 242 46
rect 274 45 275 48
rect 279 46 280 47
rect 282 46 283 48
rect 280 45 281 46
rect 277 40 282 41
rect 285 40 287 41
rect 0 35 4 39
rect 35 35 39 39
rect 238 35 242 39
rect 2 33 3 35
rect 83 33 84 35
rect 100 33 101 35
rect 2 28 3 30
rect 67 28 71 30
rect 73 28 74 29
rect 238 28 242 32
rect 257 31 258 33
rect 40 25 42 28
rect 74 27 76 28
rect 76 26 77 27
rect 83 25 84 27
rect 257 26 258 28
rect 0 21 4 25
rect 33 24 42 25
rect 25 23 42 24
rect 25 21 39 23
rect 25 20 37 21
rect 31 18 32 20
rect 37 18 38 19
rect 35 16 37 18
rect 10 13 11 14
rect 26 13 27 14
rect 28 13 29 15
rect 40 13 42 23
rect 50 20 52 23
rect 238 21 242 25
rect 294 21 295 23
rect 53 16 55 20
rect 67 13 68 14
rect 91 13 92 14
rect 9 12 10 13
rect 27 12 29 13
rect 65 12 67 13
rect 92 12 93 13
rect 28 11 30 12
rect 64 11 65 12
rect 265 11 266 12
rect 281 11 282 12
rect 0 7 4 11
rect 9 10 10 11
rect 28 10 29 11
rect 92 10 93 11
rect 10 9 11 10
rect 91 9 92 10
rect 18 8 19 9
rect 75 8 76 9
rect 19 7 21 8
rect 73 7 75 8
rect 238 7 242 11
rect 264 10 265 11
rect 282 10 284 11
rect 284 9 285 10
rect 264 8 265 9
rect 265 7 266 8
rect 21 6 22 7
rect 72 6 73 7
rect 273 6 274 7
rect 274 5 276 6
rect 276 4 277 5
use buf_1of2 b0
timestamp 906617853
transform 1 0 -300 0 1 -103
box 300 103 402 287
use router_generated_wiring gen_wiring
timestamp 976159201
transform 1 0 0 0 1 0
box -7 -143 242 81
use buf_1of2 b1
timestamp 906617853
transform 1 0 -45 0 1 -105
box 300 103 402 287
<< end >>
