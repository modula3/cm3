magic
tech scmos
timestamp 1065832382
<< ntransistor >>
rect 5 4 7 20
rect 10 4 12 20
<< ptransistor >>
rect 5 32 7 58
rect 13 32 15 58
<< ndiffusion >>
rect 0 13 5 20
rect 4 4 5 13
rect 7 4 10 20
rect 12 16 13 20
rect 12 4 15 16
<< pdiffusion >>
rect 4 49 5 58
rect 2 32 5 49
rect 7 36 13 58
rect 7 32 8 36
rect 12 32 13 36
rect 15 49 16 58
rect 15 32 18 49
<< ndcontact >>
rect 0 4 4 13
rect 13 16 17 20
<< pdcontact >>
rect 0 49 4 58
rect 8 32 12 36
rect 16 49 20 58
<< polysilicon >>
rect 5 58 7 61
rect 13 58 15 61
rect 5 29 7 32
rect 0 25 7 29
rect 13 29 15 32
rect 13 27 20 29
rect 5 20 7 25
rect 10 25 20 27
rect 10 20 12 25
rect 5 1 7 4
rect 10 1 12 4
<< genericcontact >>
rect 1 26 3 28
rect 17 26 19 28
<< metal1 >>
rect -2 60 22 65
rect 0 58 4 60
rect 16 58 20 60
rect 9 29 12 32
rect 0 24 4 29
rect 8 24 12 29
rect 16 24 20 29
rect 9 20 12 24
rect 9 17 13 20
rect 0 1 4 4
rect -2 -3 22 1
<< labels >>
rlabel metal1 2 27 2 27 1 i0
rlabel metal1 18 27 18 27 1 i1
rlabel metal1 10 27 10 27 1 o0
rlabel space -2 -5 22 67 1 _
rlabel metal1 0 -1 0 -1 2 GND!
rlabel metal1 0 63 0 63 3 Vdd!
rlabel ndiffusion 4 4 15 17 1 nwidth_north@
rlabel pdiffusion 4 35 16 58 1 pwidth_south@
<< end >>
