magic
tech scmos
timestamp 975640201
<< metal1 >>
rect 0 0 3 3
<< labels >>
rlabel metal1 1 1 1 1 1 x
<< end >>
