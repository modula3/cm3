magic
tech scmos
timestamp 1051683898
<< metal1 >>
rect -8 40 11 43
rect -8 27 -5 40
rect 0 32 4 37
rect 8 27 11 40
rect -8 24 11 27
rect 0 8 4 13
rect 16 8 20 13
rect 0 0 4 5
rect 16 0 20 5
<< labels >>
rlabel metal1 2 2 2 2 3 x
rlabel metal1 17 2 17 2 7 x
rlabel metal1 2 10 2 10 4 y
rlabel metal1 17 10 17 10 6 y
rlabel metal1 2 34 2 34 4 y
<< end >>
