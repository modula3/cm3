magic
tech scmos
timestamp 974270785
use b b_0
array 10 0 8 0 0 4
timestamp 908305645
transform 1 0 0 0 1 0
box 0 0 4 4
<< end >>
