magic
tech scmos
timestamp 0
use router_generated_wiring gen_wiring
timestamp 976094166
transform 1 0 0 0 1 0
box 0 -59 242 39
<< metal1 >>
rect 154 -63 157 -56
rect 147 -63 150 -56
rect 140 -63 143 -56
rect 133 -63 136 -56
rect 126 -63 129 -56
rect 224 0 231 3
rect 35 0 42 3
rect 0 0 7 3
rect 224 7 231 10
rect 35 7 42 10
rect 0 7 7 10
rect 224 14 231 17
rect 35 14 42 17
rect 0 14 7 17
rect 224 21 231 24
rect 35 21 42 24
rect 0 21 7 24
rect 224 28 231 31
rect 35 28 42 31
rect 0 28 7 31
<< labels >>
rlabel metal1 227 2 227 2 1 x5
rlabel metal1 227 9 227 9 5 x4
rlabel metal1 227 16 227 16 5 x3
rlabel metal1 227 23 227 23 5 x2
rlabel metal1 227 30 227 30 5 x1
rlabel metal1 155 -59 155 -59 7 x5
rlabel metal1 148 -59 148 -59 3 x4
rlabel metal1 141 -59 141 -59 3 x3
rlabel metal1 134 -59 134 -59 3 x2
rlabel metal1 127 -59 127 -59 3 x1
rlabel metal1 38 29 38 29 5 x5
rlabel metal1 38 22 38 22 1 x4
rlabel metal1 38 15 38 15 1 x3
rlabel metal1 38 8 38 8 1 x2
rlabel metal1 38 1 38 1 1 x1
rlabel metal1 3 29 3 29 5 x5
rlabel metal1 3 22 3 22 1 x4
rlabel metal1 3 15 3 15 1 x3
rlabel metal1 3 8 3 8 1 x2
rlabel metal1 3 1 3 1 1 x1
<< end >>
