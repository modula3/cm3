magic
tech scmos
timestamp 1051739388
<< metal1 >>
rect -3575 3327 -3571 3332
rect -106 2924 -102 2929
rect 1894 2865 1898 2870
rect -4889 2084 -4885 2089
rect -1977 2001 -1973 2006
rect 4025 1764 4029 1769
rect 1586 1385 1590 1390
rect -1551 687 -1547 692
rect 4842 438 4846 443
rect -2024 414 -2020 419
rect 0 0 4 5
rect 1006 -12 1010 -7
rect -3847 -225 -3843 -220
rect -154 -947 -150 -942
rect 1658 -1065 1662 -1060
rect 1101 -1172 1105 -1167
rect -1882 -1314 -1878 -1309
rect -3776 -2403 -3772 -2398
rect -982 -2438 -978 -2433
rect 2415 -2758 2419 -2753
rect -3433 -2829 -3429 -2824
rect 1326 -2912 1330 -2907
<< labels >>
rlabel metal1 1 3 1 3 3 x
rlabel metal1 -2023 417 -2023 417 3 x
rlabel metal1 1895 2868 1895 2868 3 x
rlabel metal1 -1881 -1311 -1881 -1311 3 x
rlabel metal1 -4888 2087 -4888 2087 3 x
rlabel metal1 1587 1388 1587 1388 3 x
rlabel metal1 -1976 2004 -1976 2004 3 x
rlabel metal1 4843 441 4843 441 3 x
rlabel metal1 2416 -2755 2416 -2755 3 x
rlabel metal1 -3432 -2826 -3432 -2826 3 x
rlabel metal1 1102 -1169 1102 -1169 3 x
rlabel metal1 -3846 -222 -3846 -222 3 x
rlabel metal1 1007 -9 1007 -9 3 x
rlabel metal1 -105 2927 -105 2927 3 x
rlabel metal1 -3574 3330 -3574 3330 3 x
rlabel metal1 4026 1767 4026 1767 3 x
rlabel metal1 1659 -1062 1659 -1062 3 x
rlabel metal1 -1550 690 -1550 690 3 x
rlabel metal1 -981 -2435 -981 -2435 3 x
rlabel metal1 -3775 -2400 -3775 -2400 3 x
rlabel metal1 -153 -944 -153 -944 3 x
rlabel metal1 1327 -2909 1327 -2909 3 x
<< end >>
