magic
tech scmos
timestamp 956777167
<< labels >>
rlabel space -11 -8 12 16 4 whole_cell
<< end >>
