magic
tech scmos
timestamp 1036525394
<< metal1 >>
rect 0 24 8 27
rect -8 16 16 19
rect -8 -5 -5 16
rect 0 8 8 11
rect 0 0 8 3
rect 13 -5 16 16
rect 32 0 40 3
rect -8 -8 16 -5
<< metal2 >>
rect -8 -8 16 3
use test4_sub s
timestamp 1036525394
transform 1 0 56 0 1 0
box 0 0 8 3
<< labels >>
rlabel metal1 5 9 5 9 4 y
rlabel metal1 35 2 35 2 8 y
rlabel metal1 3 1 3 1 2 x
rlabel metal1 3 25 3 25 2 x
<< end >>
