magic
tech scmos
timestamp 1035933170
<< metal1 >>
rect 0 16 7 20
rect 24 16 31 20
rect 40 16 47 20
rect 0 0 7 4
rect 24 0 31 4
rect 40 0 47 4
rect 0 -6 47 -3
<< metal2 >>
rect 0 -6 47 14
<< labels >>
rlabel metal1 4 2 4 2 1 y
rlabel metal1 4 18 4 18 2 z
rlabel metal1 28 18 28 18 1 x
rlabel metal1 27 2 27 2 1 x
rlabel metal1 43 18 43 18 1 y
rlabel metal1 43 2 43 2 8 z
<< end >>
