magic
tech scmos
timestamp 973571252
use b b_0
array 0 3 10 0 0 8
timestamp 908305645
transform -1 0 32 0 -1 8
box 0 0 4 4
<< end >>
