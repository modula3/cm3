magic
tech scmos
timestamp 1065832382
<< ntransistor >>
rect 5 4 7 20
<< ptransistor >>
rect 5 32 7 58
<< ndiffusion >>
rect 2 13 5 20
rect 4 4 5 13
rect 7 16 8 20
rect 7 4 10 16
<< pdiffusion >>
rect 4 49 5 58
rect 2 32 5 49
rect 7 36 10 58
rect 7 32 8 36
<< ndcontact >>
rect 0 4 4 13
rect 8 16 12 20
<< pdcontact >>
rect 0 49 4 58
rect 8 32 12 36
<< polysilicon >>
rect 5 58 7 61
rect 5 29 7 32
rect 0 25 7 29
rect 5 20 7 25
rect 5 1 7 4
<< genericcontact >>
rect 1 26 3 28
<< metal1 >>
rect -2 60 14 65
rect 0 58 4 60
rect 9 29 12 32
rect 0 24 4 29
rect 8 24 12 29
rect 9 20 12 24
rect 0 1 4 4
rect -2 -3 14 1
<< labels >>
rlabel metal1 -1 -1 -1 -1 2 GND!
rlabel metal1 0 63 0 63 4 Vdd!
rlabel metal1 2 27 2 27 1 i0
rlabel metal1 10 27 10 27 1 o0
rlabel space -2 -5 14 67 1 _
rlabel pdiffusion 4 35 10 58 1 pwidth_south@
rlabel ndiffusion 4 4 10 17 1 nwidth_north@
<< end >>
