magic
tech scmos
timestamp 908305645
<< polysilicon >>
rect 0 0 2 2
<< metal1 >>
rect 0 0 4 4
<< end >>
